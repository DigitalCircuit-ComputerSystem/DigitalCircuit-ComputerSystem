module cpu(
	input rst;
	input clk;
	input[31:0] data_rom_i;  //指令文件
	output[31:0] addr_rom_o;
)

wire pc;

wire[5:0]alu;  
wire [31:0]seq_pc;
wire is_jmp;
wire [31:0] jmp_pc;
wire [31:0] src1;     //值
wire [31:0] src2;
wire [31:0] dest;
wire [33:0] src1_type;  //高两位为类型 ，00：无， 01：寄存器，此时type低5位为寄存器号， 10：内存，此时type低32位为内存地址  11：常数
wire [33:0] src2_type;
wire [33:0] dest_type;
wire [31:0] src1_data;
wire [31:0] src2_data;

wire [31:0] read_data1;
wire [31:0] read_data2;
wire [31:0] write_data;
wire [4:0] write_reg;
wire [4:0] read_reg1;  //读的寄存器的地址
wire [4:0] read_reg2;
wire wr_en;  //写寄存器使能端
wire read_en1;  //读寄存器使能端
wire read_en2;

fetch_pc fetch_pc0 (.rst(rst), .clk(clk), .pc_i(pc), .is_jmp(is_jmp), .jmp_pc(jmp_pc), .pc_o(pc));  //取指令以及更新pc

decode decode0 (.ins(data_rom_i), .PC(pc), .reg1_data(read_data1), .reg2_data(read_data2), .wraddr(write_reg),
	.reg1_addr(read_reg1), .reg2_addr(read_reg2), .jmp_addr(jmp_pc), .wreg(wr_en), .is_jmp(is_jmp),
	.reg1_read(read_en1), .reg2_read(read_en2), .wdata(write_data);

regs regs0 (.clk(clk), .write_data(write_data), .write_reg(write_reg), .write_en(wr_en), .read_reg1(read_reg1),
	.read_en1(read_en1), .read_reg2(read_reg2), .read_en2(read_en2), .read_data1_o(read_data1), .read_data2_o(read_data2));

